-- This file is part of the Omega CPU Core
-- Copyright 2015 - 2016 Joseph Shetaye

-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU Lesser General Public License as
-- published by the Free Software Foundation, either version 3 of the
-- License, or (at your option) any later version.

-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.

-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.

library IEEE;
use IEEE.std_logic_1164.all;
use work.constants.all;
use IEEE.Numeric_std.all;

entity MemoryController is

  port (
    CLK         : in  std_logic;
    Address     : in  word;
    Enable      : in  std_logic;
    ToWrite     : in  word;
    FromRead    : out word;
    Instruction : in  word;
    Reset       : in  std_logic;
    Done        : out std_logic;
	 SRAM_addr     : out std_logic_vector(20 downto 0);
    SRAM_OE       : out std_logic;
    SRAM_CE       : out std_logic;
    SRAM_WE       : out std_logic;
    SRAM_data     : inout  std_logic_vector(7 downto 0);
	 Status_Debug  : out std_logic_vector(7 downto 0)
	 );
  
end MemoryController;

architecture Behavioral of MemoryController is

 constant LoadByteUnsigned : Operator := "000";
 constant LoadByteSigned : Operator := "001";
 constant LoadHalfWordUnsigned : Operator := "010";
 constant LoadHalfWordSigned : Operator := "011";
 constant LoadWord : Operator := "100";
 constant StoreByte : Operator := "101";
 constant StoreHalfWord : Operator := "110";
 constant StoreWord : Operator := "111";
 
 -- Put boot image here
 --constant BootImage : MemoryArray := ();
 
 constant BootImage : MemoryArray := ("01000011","00000000","00100000","00100100","00000000","00000000","01000000","00100100","00001000","00000000","01000010","01010100",
"00000000","00000000","01000010","00100100","00001000","00000000","01000010","01010100","00000000","00000000","01000010","00100100","00001000","00000000","01000010","01010100",
"01000100","00000000","01000010","00100100","00000000","00000000","00100010","10011100","00000000","00000000","00100000","00100000","00000000","00000000","00100010","10010000",
"00000000","00000000","00100001","10110100","00000000","00000000","01100000","00100000","00000001","00000000","01100011","00100100","11101000","00000011","10000011","01100100",
"11111110","11111111","10011111","11010000","11110000","11111111","11111111","11001011","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000",
"00000000","00000000","00000000");

 signal FromRead_S : Word := (others => '0');
 signal NeedsInit : std_logic := '1';
 signal BootImageIndex : Integer := 0;
 signal Done_s : std_logic := '0';
 signal SRAM_addr_s : std_logic_vector(20 downto 0) := (others => '0');
 signal SRAM_data_s : std_logic_vector(7 downto 0); --:= (others => 'Z');
 signal SRAM_datain_s : std_logic_vector(7 downto 0);
 signal SRAM_bootloaderData_s : std_logic_vector(7 downto 0);
 signal SRAM_OE_s : std_logic := '1';
 signal SRAM_WE_s : std_logic := '1';
 signal SRAM_CE_s : std_logic := '1';
 signal AddressOffset : integer := 0;
 --signal Status_Debug_s : std_logic_vector(7 downto 0) := (others => '0');
begin  -- Behavioral

  SRAM_addr <= SRAM_addr_s;
  --SRAM_data <= SRAM_bootloaderData_s when SRAM_OE_s = '1' else (others => 'Z');
  SRAM_datain_s <= SRAM_data when SRAM_OE_s = '0' else (others => '0');
  SRAM_OE <= SRAM_OE_s;
  SRAM_WE <= SRAM_WE_s;
  SRAM_CE <= '0';
    FromRead <= FromRead_S;
	 Done <= Done_s;
	 --Status_Debug <= Status_Debug_S;
	 
  process (CLK)
  begin
	if SRAM_OE_s = '0' then
		SRAM_data <= (others => 'Z');
   elsif NeedsInit = '1' then
		SRAM_data <= SRAM_bootloaderData_s;
	else
		SRAM_data <= SRAM_data_s;
	end if;
  end process;
  
  process (CLK)--(Enable, Instruction, Address, Reset)
	-- Removed procedure initialize
	  variable current_operator : std_logic_vector(2 downto 0);
  begin  -- process
  if rising_edge(CLK) then
    if NeedsInit = '1' then
	   if BootImageIndex = BootImage'Length then
			SRAM_we_s <= '1';
			NeedsInit <= '0';
			SRAM_oe_s <= '1';
		else
			SRAM_bootloaderData_s <= BootImage(BootImageIndex);
			SRAM_addr_s <= std_logic_vector(to_unsigned(BootImageIndex,21));
		   SRAM_we_s <= '0';
			BootImageIndex <= BootImageIndex + 1;
		end if;
    elsif Enable = '1' then
	 current_operator := GetOperator(Instruction);
    case current_operator is
      when LoadByteUnsigned =>
		  if SRAM_oe_s = '1' then
				SRAM_addr_s <= Address(20 downto 0);
				SRAM_oe_s <= '0';
				Done_s <= '0';
			else
				FromRead_S <= "000000000000000000000000" & SRAM_datain_s;
				SRAM_oe_s <= '1';
				Done_s <= '1';
			end if;
      when LoadByteSigned =>
		  if SRAM_oe_s = '1' then
				SRAM_addr_s <= Address(20 downto 0);
				SRAM_oe_s <= '0';
				Done_s <= '0';
			else
				FromRead_S <= std_logic_vector(resize(signed(SRAM_datain_s),32));
				SRAM_oe_s <= '1';
				Done_s <= '1';
			end if;
      when LoadHalfWordUnsigned =>
			if SRAM_oe_s = '1' then
				SRAM_addr_s <= Address(20 downto 0);
				SRAM_oe_s <= '0';
				AddressOffset <= 0;
				Done_s <= '0';
		   elsif AddressOffset < 1 then
				SRAM_addr_s <= std_logic_vector(unsigned(Address(20 downto 0)) + to_unsigned(AddressOffset + 1,20));
				AddressOffset <= AddressOffset + 1;
				FromRead_S(8*AddressOffset+7 downto 8*AddressOffset) <= SRAM_datain_s;
			else
				FromRead_S(8*AddressOffset+7 downto 8*AddressOffset) <= SRAM_datain_s;
				FromRead_S(31 downto 16) <= (others => '0');
				AddressOffset <= 0;
				SRAM_oe_s <= '1';
				Done_s <= '1';
			end if;
      when LoadHalfWordSigned =>
			if SRAM_oe_s = '1' then
				SRAM_addr_s <= Address(20 downto 0);
				SRAM_oe_s <= '0';
				AddressOffset <= 0;
				Done_s <= '0';
		   elsif AddressOffset < 1 then
				SRAM_addr_s <= std_logic_vector(unsigned(Address(20 downto 0)) + to_unsigned(AddressOffset + 1,20));
				AddressOffset <= AddressOffset + 1;
				FromRead_S(8*AddressOffset+7 downto 8*AddressOffset) <= SRAM_datain_s;
			else
				FromRead_S(8*AddressOffset+7 downto 8*AddressOffset) <= SRAM_datain_s;
				if SRAM_datain_s(7) = '1' then
				   FromRead_S(31 downto 16) <= "1111111111111111";
				else
				   FromRead_S(31 downto 16) <= "0000000000000000";
				end if;
				AddressOffset <= 0;
				SRAM_oe_s <= '1';
				Done_s <= '1';
			end if;
      when LoadWord =>
			if SRAM_oe_s = '1' then
				SRAM_addr_s <= Address(20 downto 0);
				SRAM_oe_s <= '0';
				AddressOffset <= 0;
				Done_s <= '0';
		   elsif AddressOffset < 3 then
				SRAM_addr_s <= std_logic_vector(unsigned(Address(20 downto 0)) + to_unsigned(AddressOffset+1,20));
				FromRead_S(8*AddressOffset+7 downto 8*AddressOffset) <= SRAM_datain_s;
				AddressOffset <= AddressOffset + 1;
			else
				FromRead_S(8*AddressOffset+7 downto 8*AddressOffset) <= SRAM_datain_s;
				AddressOffset <= 0;
				SRAM_oe_s <= '1';
				Done_s <= '1';
				--Status_Debug_S <= Address(9 downto 2) xor "11111111";
			end if;
      when StoreByte =>
			SRAM_oe_s <= '1';
			if SRAM_we_s = '1' then
				SRAM_addr_s <= Address(20 downto 0);
				SRAM_data_s <= ToWrite(7 downto 0);
				SRAM_we_s <= '0';
			else
				SRAM_we_s <= '1';
				Done_s <= '1';
			end if;
 --      Memory(to_integer(unsigned(Address))) <= ToWrite(7 downto 0);
      when StoreHalfWord =>
			SRAM_oe_s <= '1';
			if SRAM_we_s = '1' then
				SRAM_addr_s <= Address(20 downto 0);
				SRAM_data_s <= ToWrite(7 downto 0);
				SRAM_we_s <= '0';
				Done_s <= '0';
			elsif AddressOffset < 1 then
				SRAM_addr_s <= std_logic_vector(unsigned(Address(20 downto 0)) + to_unsigned(AddressOffset+1,20));
				SRAM_data_s <= ToWrite(8*AddressOffset+7 downto 8*AddressOffset);
				AddressOffset <= AddressOffset + 1;
			else
				AddressOffset <= 0;
				SRAM_we_s <= '1';
				Done_s <= '1';
			end if;
--        Memory(to_integer(unsigned(Address))) <= ToWrite(7 downto 0);
--        Memory(to_integer(unsigned(Address)) + 1) <= ToWrite(15 downto 8);
      when StoreWord =>
			SRAM_oe_s <= '1';
			if SRAM_we_s = '1' then
				SRAM_addr_s <= Address(20 downto 0);
				SRAM_data_s <= ToWrite(7 downto 0);
				SRAM_we_s <= '0';
				Done_s <= '0';
			elsif AddressOffset < 3 then
				SRAM_addr_s <= std_logic_vector(unsigned(Address(20 downto 0)) + to_unsigned(AddressOffset+1,20));
				SRAM_data_s <= ToWrite(8*AddressOffset+7 downto 8*AddressOffset);
				AddressOffset <= AddressOffset + 1;
			else
				AddressOffset <= 0;
				SRAM_we_s <= '1';
				Done_s <= '1';
			end if;
--        Memory(to_integer(unsigned(Address))) <= ToWrite(7 downto 0);
--        Memory(to_integer(unsigned(Address)) + 1) <= ToWrite(15 downto 8);
--        Memory(to_integer(unsigned(Address)) + 2) <= ToWrite(23 downto 16);
--        Memory(to_integer(unsigned(Address)) + 3) <= ToWrite(31 downto 24);
      when others => null;
    end case;
  else
    SRAM_oe_s <= '1';
	 SRAM_we_s <= '1';
    Done_s <= '0';
  end if;
  end if;
  end process;

end Behavioral;
