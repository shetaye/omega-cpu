 -- outputTest (absolute jump)
 --constant BootImage : MemoryArray := ("01000001","00000000","00100000","00100100","00000000","00000000","00100001","10110100","00000001","00000000","00000000","11000100","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000");
 -- outputTest (relative jump)
 --constant BootImage : MemoryArray := ("01000001","00000000","00100000","00100100","00000000","00000000","00100001","10110100","11111111","11111111","11111111","11001011","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000");
 -- ROT13
 --constant BootImage : MemoryArray := ("00000000","00000000","10000001","10100100","01000001","00000000","00100100","01110100","00001010","00000000","00100000","11011000","01011011","00000000","00100100","01110100","00001001","00000000","00100000","11011000","01100001","00000000","00100100","01110100","00000110","00000000","00100000","11011000","01111011","00000000","00100100","01110100","00001100","00000000","00100000","11011000","00000011","00000000","00000000","11001000","00000000","00000000","10000001","10110100","11110101","11111111","11111111","11001011","11111110","11111111","11111111","11001011","10111111","11111111","10000100","00100100","00001101","00000000","10000100","00100100","00011010","00000000","00100100","01110100","00000010","00000000","00100000","11011000","11100110","11111111","10000100","00100100","01000001","00000000","10000100","00100100","11110111","11111111","11111111","11001011","10011111","11111111","10000100","00100100","00001101","00000000","10000100","00100100","00011010","00000000","00100100","01110100","00000010","00000000","00100000","11011000","11100110","11111111","10000100","00100100","01100001","00000000","10000100","00100100","11110000","11111111","11111111","11001011","00000000","00000000","00000000");--(others => (others => '0'));
 -- Divide Test
 --constant BootImage : MemoryArray := ("10100000","00001111","01100000","00100111","00000001","00000000","00000000","11001000","00000000","00000000","10000001","10100100","00000000","00000000","10100001","10100100","01000000","00101001","10000100","00111000","00000000","00000000","10000001","10110100","00000000","00000000","10100001","10110100","11111011","11111111","11111111","11001011", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000");
 -- Output A Test 
 --constant BootImage : MemoryArray := ("01000001","00000000","00100000","00100100","00000000","00000000","00100001","10110100","11111111","11111111","11111111","11001011","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000");
 -- Echo
 --constant BootImage : MemoryArray := ("00000000","00000000","00100001","10100100","00000000","00000000","00100001","10110100","11111110","11111111","11111111","11001011","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000");
 -- Echo A-Z
 --constant BootImage : MemoryArray := ("01000000","00000000","01000000","00100100","00000001","00000000","01000010","00100100","01011011","00000000","01100010","00101100","00000110","00000000","01100000","11010000","00000001","00000000","10000100","00100100","01010000","11000011","10100100","00101100","11111110","11111111","10111111","11011000","00000000","00000000","01000001","10110100","11111001","11111111","11111111","11001011","01000000","00000000","01000000","00100100","11111010","11111111","11111111","11001011","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000");
 -- Output B Test
 --constant BootImage :  MemoryArray := ("01000010","00000000","00100000","00100100","00000011","00000000","00000000","11001000","00000000","00000000","00100001","10110100","11111110","11111111","11111111","11001011","11101000","00000011","10000000","00100100","00000000","00000000","10100000","00100100","00000001","00000000","10100101","00100100","00000000","00101000","11000100","01100000","11111110","11111111","11011111","11010000","11111001","11111111","11111111","11001011","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000");
 -- Calculator Demo
 constant BootImage : MemoryArray := ("01010011","01111001","01101110","01110100","01100001","01111000","00100000","01100101","01110010","01110010","01101111","01110010","00001010","00000000","00000000","00000000","01000100","01101001","01110110","01101001","01100100","01100101","00100000","01100010","01111001","00100000","01111010","01100101","01110010","01101111","00001010","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000110","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000111","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00001000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00010000","00000000","00000000","00000000","00010001","00000000","00000000","00000000","00010010","00000000","00000000","00000000","00010011","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00100100","00000000","00001000","00100101","00000000","00000000","00101000","10010001","00001100","00000000","00100000","11010001","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101000","00000000","01001010","00100101","00000000","00000000","01100000","10100101","00000000","00000000","01001011","10011101","00000000","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00100000","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000001","00000000","00101001","00100101","00001000","00000000","00101001","01010101","01011000","00000000","00101001","00100101","00000100","00000000","00001000","00110101","00000000","01000000","00101001","00100001","00000000","00000000","00001001","11000000","00000101","00000000","00000000","11001000","00000101","00000000","00000000","11001000","11001100","00000000","00000000","11001000","00011101","00000001","00000000","11001000","00101011","00000001","00000000","11001000","01111010","00000001","00000000","11001000","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00101000","00000000","00001000","00100101","00000000","00000000","00101000","10010001","00110000","00000000","01001001","01100101","00100100","00000000","01000000","11010001","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00100000","00000000","01001010","00100101","00000011","00000000","01100000","00100101","00000000","00000000","01001011","10011101","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00110000","00000000","01001010","00100101","00000000","00000000","01100000","00100101","00000000","00000000","01001011","10011101","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101000","00000000","01001010","00100101","00000000","00000000","01001010","10010001","00000000","00000000","01100000","00100101","00001000","00000000","01101011","01010101","00000000","00000000","01101011","00100101","00001000","00000000","01101011","01010101","00000000","00000000","01101011","00100101","00001000","00000000","01101011","01010101","00101100","00000000","01101011","00100101","00000000","00000000","01101010","10011101","01001101","00000001","00000000","11001000","00110001","00000000","01001001","01110101","11111111","11111111","10001001","00110101","11000110","11111111","01100010","01110101","00000000","01011000","01001010","00000001","00110110","00000000","01000000","11010001","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00100000","00000000","01001010","00100101","00000000","00000000","01101010","10010001","00000010","00000000","01100000","00100101","00000000","00000000","01001011","10011101","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101000","00000000","01001010","00100101","00000000","00000000","01101010","10010001","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00110000","00000000","01001010","00100101","00110000","00000000","01101011","00101101","00000000","00000000","01001011","10011101","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101000","00000000","01001010","00100101","00000000","00000000","01001010","10010001","00000000","00000000","01100000","00100101","00001000","00000000","01101011","01010101","00000000","00000000","01101011","00100101","00001000","00000000","01101011","01010101","00000000","00000000","01101011","00100101","00001000","00000000","01101011","01010101","00101100","00000000","01101011","00100101","00000000","00000000","01101010","10011101","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101000","00000000","01001010","00100101","00000000","00000000","01100001","10100101","00000000","00000000","01001011","10011101","00010011","00000001","00000000","11001000","00101011","00000000","01001001","01100101","00101101","00000000","01101001","01100101","00000000","01011000","01001010","00000001","00101010","00000000","01101001","01100101","00000000","01011000","01001010","00000001","00101111","00000000","01101001","01100101","00000000","01011000","01001010","00000001","00101000","00000000","01101001","01100101","00000000","01011000","01001010","00000001","00101001","00000000","01101001","01100101","00000000","01011000","01001010","00000001","00100100","00000000","01000000","11010001","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00100000","00000000","01001010","00100101","00000100","00000000","01100000","00100101","00000000","00000000","01001011","10011101","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101000","00000000","01001010","00100101","00000000","00000000","01001010","10010001","00000000","00000000","01100000","00100101","00001000","00000000","01101011","01010101","00000000","00000000","01101011","00100101","00001000","00000000","01101011","01010101","00000000","00000000","01101011","00100101","00001000","00000000","01101011","01010101","00101100","00000000","01101011","00100101","00000000","00000000","01101010","10011101","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101000","00000000","01001010","00100101","00000000","00000000","01100001","10100101","00000000","00000000","01001011","10011101","11100100","00000000","00000000","11001000","00100000","00000000","01001001","01100101","00001001","00000000","01101001","01100101","00000000","01011000","01001010","00000001","00010100","00000000","01000000","11010001","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00100000","00000000","01001010","00100101","00000001","00000000","01100000","00100101","00000000","00000000","01001011","10011101","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101000","00000000","01001010","00100101","00000000","00000000","01100001","10100101","00000000","00000000","01001011","10011101","11001101","00000000","00000000","11001000","00001010","00000000","01001001","01100101","00001101","00000000","01000000","11010001","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00100100","00000000","01001010","00100101","00000001","00000000","01100000","00100101","00000000","00000000","01001011","10011101","00001000","00000000","01000000","00100101","00000000","00000000","10001010","10011100","00000000","00000000","00011101","11000000","00000000","00000000","00011101","11000000","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00100100","00000000","01001010","00100101","00000001","00000000","01100000","00100101","00000000","00000000","01001011","10011101","00000111","00000000","01000000","00100101","00000000","00000000","10001010","10011100","00000000","00000000","00011101","11000000","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00101000","00000000","00101001","00100101","00000000","00000000","00101001","10010001","00110000","00000000","01001001","01110101","11111111","11111111","10001001","00110101","11000111","11111111","01101100","01110101","00000000","01011000","01001010","00000001","00111000","00000000","01000000","11011001","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00110000","00000000","01001010","00100101","00000000","00000000","01101010","10010001","00001010","00000000","01101011","00110101","00000000","00000000","01001011","10011101","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101000","00000000","01001010","00100101","00000000","00000000","01001010","10010001","00110000","00000000","01001010","00101101","00000000","00000000","01100000","00100101","00001000","00000000","01101011","01010101","00000000","00000000","01101011","00100101","00001000","00000000","01101011","01010101","00000000","00000000","01101011","00100101","00001000","00000000","01101011","01010101","00110000","00000000","01101011","00100101","00000000","00000000","10001011","10010001","00000000","01100000","01001010","00100001","00000000","00000000","01101010","10011101","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101000","00000000","01001010","00100101","00000000","00000000","01001010","10010001","00000000","00000000","01100000","00100101","00001000","00000000","01101011","01010101","00000000","00000000","01101011","00100101","00001000","00000000","01101011","01010101","00000000","00000000","01101011","00100101","00001000","00000000","01101011","01010101","00101100","00000000","01101011","00100101","00000000","00000000","01101010","10011101","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101000","00000000","01001010","00100101","00000000","00000000","01100001","10100101","00000000","00000000","01001011","10011101","01101110","00000000","00000000","11001000","00000000","00000000","01000000","00100101","00000000","00000000","10001010","10011100","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00110000","00000000","01001010","00100101","00000000","00000000","01001010","10010001","00000100","00000000","01100100","00100101","00000000","00000000","01101010","10011101","00000000","00000000","00011101","11000000","01100000","00000000","00000000","11001000","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00100000","00000000","01001010","00100101","00000001","00000000","01100000","00100101","00000000","00000000","01001011","10011101","00000000","00000000","01000000","00100101","00000000","00000000","10001010","10011100","00000100","00000000","01100100","00100101","00000000","00000000","01100000","10011101","00000000","00000000","00011101","11000000","01010001","00000000","00000000","11001000","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00100000","00000000","01001010","00100101","00000001","00000000","01100000","00100101","00000000","00000000","01001011","10011101","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101100","00000000","01001010","00100101","00000000","00000000","01001010","10010001","00101011","00000000","01001010","01100101","00000100","00000000","01000000","11010001","00000001","00000000","01000000","00100101","00000000","00000000","10001010","10011100","00110111","00000000","00000000","11001000","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101100","00000000","01001010","00100101","00000000","00000000","01001010","10010001","00101101","00000000","01001010","01100101","00000100","00000000","01000000","11010001","00000010","00000000","01000000","00100101","00000000","00000000","10001010","10011100","00101010","00000000","00000000","11001000","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101100","00000000","01001010","00100101","00000000","00000000","01001010","10010001","00101111","00000000","01001010","01100101","00000100","00000000","01000000","11010001","00000100","00000000","01000000","00100101","00000000","00000000","10001010","10011100","00011101","00000000","00000000","11001000","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101100","00000000","01001010","00100101","00000000","00000000","01001010","10010001","00101010","00000000","01001010","01100101","00000100","00000000","01000000","11010001","00000011","00000000","01000000","00100101","00000000","00000000","10001010","10011100","00010000","00000000","00000000","11001000","00000000","00000000","01000000","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00000000","00000000","01001010","00100101","00001000","00000000","01001010","01010101","00101100","00000000","01001010","00100101","00000000","00000000","01001010","10010001","00101000","00000000","01001010","01100101","00000100","00000000","01000000","11010001","00000101","00000000","01000000","00100101","00000000","00000000","10001010","10011100","00000011","00000000","00000000","11001000","00000110","00000000","01000000","00100101","00000000","00000000","10001010","10011100","00000100","00000000","01000100","00100101","00000000","00000000","01000000","10011101","00000000","00000000","00011101","11000000","00000001","00000000","00000000","11001000","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00100000","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000001","00000000","00001000","01100101","01100110","11111110","00011111","11010001","00000000","00000000","00011101","11000000","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10111100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000000","01000000","10100000","00100011","00000001","00000000","10111101","00101111","00000000","00000000","10100000","10011111","00000001","00000000","10111101","00101111","00000000","00000000","10100000","10011111","00000000","00000000","00011101","11000000","00000100","00000000","10111101","00101111","00000000","00000000","10100100","10011111","00000100","00000000","10111101","00101111","00000000","00000000","10100101","10011111","00000000","00000000","00011101","11000000","00000000","00000000","00011101","10010001","00000000","00000000","00000100","10011101","00000100","00000000","10111101","00100111","00000000","00000000","00011101","10010001","00000000","00000000","00000101","10011101","00000100","00000000","10111101","00100111","00000000","00000000","00011101","11000000","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00100100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00000000","00000000","00000000","10100101","00001010","00000000","00001000","01100101","11111110","11111111","00011111","11011001","00000000","00000000","00011101","11000000","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00100000","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10111100","00000000","00001000","00100101","00000000","00000000","00011101","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00100100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000000","00000000","00101000","10010001","00010100","00000000","00100000","11010001","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10001000","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","11111001","11111101","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10110000","00000000","00001000","00100101","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10001000","00000000","00101001","00100101","00000000","00000000","00101001","10010001","00000000","00000000","00001001","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10110100","00000000","00001000","00100101","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10001000","00000000","00101001","00100101","00000100","00000000","00101001","00100101","00000000","00000000","00101001","10010001","00000000","00000000","00001001","10011101","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10111000","00000000","00101001","00100101","00000000","11101000","00000000","00100001","00000100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000000","00000000","00101000","10011101","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10111000","00000000","00101001","00100101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00001001","00000000","00001000","00100101","00001000","00000000","00001000","01010101","11101100","00000000","00001000","00100101","00000000","00000000","00101001","10010001","00000100","00000000","00101001","00110101","00000000","01001000","00001000","00100001","00000000","00000000","00001000","11001100","00010010","00000000","00000000","11001000","01010101","00000010","00000000","11001000","10100000","00000000","00000000","11001000","00010111","00000001","00000000","11001000","10011110","00000000","00000000","11001000","11001110","00000010","00000000","11001000","00101001","00000001","00000000","11001000","10001000","00000010","00000000","11001000","11001110","00000001","00000000","11001000","11001010","00000010","00000000","11001000","10011000","00000000","00000000","11001000","10010111","00000000","00000000","11001000","10010110","00000000","00000000","11001000","10010101","00000000","00000000","11001000","11000101","00000010","00000000","11001000","11100100","00000010","00000000","11001000","00001000","00000100","00000000","11001000","11001110","00000100","00000000","11001000","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10110000","00000000","00101001","00100101","00000000","00000000","00101001","10010001","00000000","00000000","01001001","01100101","00011110","00000000","01000000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10110100","00000000","00101001","00100101","00000000","00000000","00101001","10010001","00000100","00000000","00001000","00100101","00000000","00000000","00001001","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01010111","00000000","00000000","11001000","00000010","00000000","01001001","01100101","00010100","00000000","01000000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00000010","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01000010","00000000","00000000","11001000","00001000","00000000","01001001","01100101","00001011","00000000","01000000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00000011","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00110110","00000000","00000000","11001000","00000101","00000000","01001001","01100101","00010100","00000000","01000000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00000100","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00100001","00000000","00000000","11001000","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","00001010","11111111","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","11100101","11111110","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00011000","00000101","00000000","11001000","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10011100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","11010111","11111110","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000101","00000101","00000000","11001000","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10110000","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000000","00000000","00101000","01100101","00011100","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10110100","00000000","00101001","00100101","00000100","00000000","00001000","00100101","00000000","00000000","00101001","10010001","00000000","00000000","00001001","10011101","00111000","00000000","00000000","11001000","00000010","00000000","00101000","01100101","00001011","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00000010","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00101100","00000000","00000000","11001000","00000101","00000000","00101000","01100101","00001010","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00000100","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","10011011","11111110","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","01110110","11111110","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00000001","00000000","00000000","11001000","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10011100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","01101000","11111110","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","10001101","00000100","00000000","11001000","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","01000101","11111110","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01111000","00000100","00000000","11001000","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10110000","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000010","00000000","00101000","01100101","00001011","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00001010","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01111001","00000000","00000000","11001000","00000001","00000000","00101000","01100101","00001011","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00001011","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01101101","00000000","00000000","11001000","00000011","00000000","00101000","01100101","00001011","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00001100","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01100001","00000000","00000000","11001000","00000100","00000000","00101000","01100101","00001011","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00001101","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01010101","00000000","00000000","11001000","00001000","00000000","00101000","01100101","00110011","00000000","00100000","11010001","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","00000010","11111110","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10100100","00000000","00101001","00100101","00000100","00000000","00101001","00100101","00000000","00000000","00101001","10010001","00110000","00000000","00101001","00100101","00000000","00000000","00100000","10110101","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","11011001","11111101","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00001100","00000100","00000000","11001000","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","11011110","11111101","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","10111001","11111101","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","11101100","00000011","00000000","11001000","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10011100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","10101011","11111101","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10110000","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000010","00000000","00101000","01100101","00001011","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00001010","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01111011","00000010","00000000","11001000","00000001","00000000","00101000","01100101","00001011","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00001011","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01101111","00000010","00000000","11001000","00000011","00000000","00101000","01100101","00001011","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00001100","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01100011","00000010","00000000","11001000","00000100","00000000","00101000","01100101","00001011","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00001101","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01010111","00000010","00000000","11001000","00000110","00000000","00101000","01100101","00001011","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00001111","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01001011","00000010","00000000","11001000","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","01011111","11111101","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","00111010","11111101","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01101101","00000011","00000000","11001000","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10011100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","00101100","11111101","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01010001","00000011","00000000","11001000","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","00010101","11111101","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","11101000","00000000","00100001","00000100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000100","00000000","00001000","00110101","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00110100","00000000","00101001","00100101","00000000","01000000","00001001","00100001","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10100100","00000000","00101001","00100101","00000000","00000000","00101000","10011101","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","11101010","11111100","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00011000","00000011","00000000","11001000","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","11011100","11111100","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000010","00000000","10111101","00100111","00000000","11101000","00000000","00100001","00000100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000100","00000000","00001000","00110101","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00110100","00000000","00101001","00100101","00000000","01000000","00001001","00100001","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10100100","00000000","00101001","00100101","00000000","00000000","00101000","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10100100","00000000","00001000","00100101","00000100","00000000","00000000","00100101","11111111","11111111","00101000","00110101","00000000","00000000","00001001","10011101","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","10100110","11111100","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","11010100","00000010","00000000","11001000","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","10100110","11111100","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","10000001","11111100","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","10110100","00000010","00000000","11001000","00000010","00000000","10111101","00100111","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","01110111","11111100","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000010","00000000","10111101","00100111","00000000","11101000","00000000","00100001","00000100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000100","00000000","00001000","00110101","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00110100","00000000","00101001","00100101","00000000","01000000","00001001","00100001","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10100100","00000000","00101001","00100101","00000000","00000000","00101000","10011101","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","01001011","11111100","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","01111001","00000010","00000000","11001000","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10011100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","00111101","11111100","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000010","00000000","10111101","00100111","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","00101010","11111100","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","11101000","00000000","00100001","00000100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000100","00000000","00001000","00110101","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00110100","00000000","00101001","00100101","00000000","01000000","00001001","00100001","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10100100","00000000","00101001","00100101","00000000","00000000","00101000","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00000100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10100100","00000000","00101001","00100101","00000100","00000000","00101001","00100101","00000000","00000000","01001001","10010001","00000000","01010000","01001000","00110001","00000000","00000000","00101010","10011101","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","11101011","11111011","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00011001","00000010","00000000","11001000","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10011100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","11011101","11111011","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000010","00000000","10111101","00100111","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","11001010","11111011","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00000100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00100001","00000000","00000000","11011001","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","10111100","11111011","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","10010111","11111011","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","11001010","00000001","00000000","11001000","00000000","11101000","00000000","00100001","00000100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000100","00000000","00001000","00110101","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00110100","00000000","00101001","00100101","00000000","01000000","00001001","00100001","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10100100","00000000","00101001","00100101","00000000","00000000","00101000","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00000100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10100100","00000000","00101001","00100101","00000100","00000000","00101001","00100101","00000000","00000000","01001001","10010001","00000000","01000000","01001010","00111001","00000000","00000000","00101010","10011101","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","01100001","11111011","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","10001111","00000001","00000000","11001000","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10110000","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000011","00000000","00101000","01100101","00000100","00000000","01001000","01100101","00000000","01001000","00101010","00000001","01011100","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10110000","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000011","00000000","00101000","01100101","00001011","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00001100","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00101101","00000000","00000000","11001000","00000100","00000000","00101000","01100101","00001011","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00001101","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00100001","00000000","00000000","11001000","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","00110101","11111011","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","00010000","11111011","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01000011","00000001","00000000","11001000","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10011100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","00000010","11111011","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10011100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","11101100","11111010","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000010","00000000","10111101","00100111","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","11011001","11111010","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","11101000","00000000","00100001","00000100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000100","00000000","00001000","00110101","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00110100","00000000","00101001","00100101","00000000","01000000","00001001","00100001","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10100100","00000000","00101001","00100101","00000000","00000000","00101000","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00000100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10100100","00000000","00101001","00100101","00000100","00000000","00101001","00100101","00000000","00000000","01001001","10010001","00000000","01000000","01001010","00101001","00000000","00000000","00101010","10011101","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","10011010","11111010","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","11001000","00000000","00000000","11001000","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10110000","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000011","00000000","00101000","01100101","00000100","00000000","01001000","01100101","00000000","01001000","00101010","00000001","01011100","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10110000","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000011","00000000","00101000","01100101","00001011","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00001100","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01100110","11111111","11111111","11001011","00000100","00000000","00101000","01100101","00001011","00000000","00100000","11010001","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00001101","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00100001","00000000","00000000","11001000","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","01101110","11111010","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","01001001","11111010","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","01111100","00000000","00000000","11001000","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10011100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","00111011","11111010","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10000100","00000000","00001000","00100101","00000001","00000000","00100000","00100101","00000000","00000000","00001001","10011101","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10011100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","00100101","11111010","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000010","00000000","10111101","00100111","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","00010010","11111010","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000000","11101000","00000000","00100001","00000100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000100","00000000","00001000","00110101","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00110100","00000000","00101001","00100101","00000000","01000000","00001001","00100001","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10100100","00000000","00101001","00100101","00000000","00000000","00101000","10011101","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10011100","00000000","00001000","00100101","00000100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000000","00000000","00100000","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","00000000","00000000","00101001","00100101","00001000","00000000","00101001","01010101","10100100","00000000","00101001","00100101","00000100","00000000","00101001","00100101","00000000","00000000","01001001","10010001","00000000","01000000","01001010","00100001","00000000","00000000","00101010","10011101","00000000","00000000","10000000","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","00000000","00000000","10000100","00100100","00001000","00000000","10000100","01010100","10100100","00000000","10000100","00100100","00000000","00000000","10011011","10011111","00000000","00000000","10011011","00100111","00000100","00000000","01111011","00101111","00000000","00000000","10111011","10011111","00000100","00000000","01111011","00101111","00000100","00000000","10111111","00100111","11010011","11111001","11111111","11001011","00000100","00000000","01111100","00101111","00000000","00000000","10111011","10010011","00000100","00000000","01111011","00100111","00000000","00000000","10011011","10010011","00000001","00000000","00000000","11001000","00000000","00000000","00000000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","00000000","00000000","00001000","00100101","00001000","00000000","00001000","01010101","10101100","00000000","00001000","00100101","00000000","00000000","00001000","10010001","00000001","00000000","00001000","00101101","11110111","11111001","00011111","11011001");
